module decoder #(parameter SIZE = 5) (
inp_i,
out_o,
);

input [SIZE-1:0] inp_i;
output [2**SIZE-1:o] out_o;

always_comb begin
	case (inp_i)
		5'h00: out_o=32'b0000_0000_0000_0000_0000_0000_0000_0001;
		5'h01: out_o=32'b0000_0000_0000_0000_0000_0000_0000_0010;
		5'h02: out_o=32'b0000_0000_0000_0000_0000_0000_0000_0100;
		5'h03: out_o=32'b0000_0000_0000_0000_0000_0000_0000_1000;
		5'h04: out_o=32'b0000_0000_0000_0000_0000_0000_0001_0000;
		5'h05: out_o=32'b0000_0000_0000_0000_0000_0000_0010_0000;
		5'h06: out_o=32'b0000_0000_0000_0000_0000_0000_0100_0000;
		5'h07: out_o=32'b0000_0000_0000_0000_0000_0000_1000_0000;
		5'h08: out_o=32'b0000_0000_0000_0000_0000_0001_0000_0000;
		5'h09: out_o=32'b0000_0000_0000_0000_0000_0010_0000_0000;
		5'h0A: out_o=32'b0000_0000_0000_0000_0000_0100_0000_0000;
		5'h0B: out_o=32'b0000_0000_0000_0000_0000_1000_0000_0000;
		5'h0C: out_o=32'b0000_0000_0000_0000_0001_0000_0000_0000;
		5'h0D: out_o=32'b0000_0000_0000_0000_0010_0000_0000_0000;
		5'h0E: out_o=32'b0000_0000_0000_0000_0100_0000_0000_0000;
		5'h0F: out_o=32'b0000_0000_0000_0000_1000_0000_0000_0000;
		5'h10: out_o=32'b0000_0000_0000_0001_0000_0000_0000_0000;
		5'h11: out_o=32'b0000_0000_0000_0010_0000_0000_0000_0000;
		5'h12: out_o=32'b0000_0000_0000_0100_0000_0000_0000_0000;
		5'h13: out_o=32'b0000_0000_0000_1000_0000_0000_0000_0000;
		5'h14: out_o=32'b0000_0000_0001_0000_0000_0000_0000_0000;
		5'h15: out_o=32'b0000_0000_0010_0000_0000_0000_0000_0000;
		5'h16: out_o=32'b0000_0000_0100_0000_0000_0000_0000_0000;
		5'h17: out_o=32'b0000_0000_1000_0000_0000_0000_0000_0000;
		5'h18: out_o=32'b0000_0001_0000_0000_0000_0000_0000_0000;
		5'h19: out_o=32'b0000_0010_0000_0000_0000_0000_0000_0000;
		5'h1A: out_o=32'b0000_0100_0000_0000_0000_0000_0000_0000;
		5'h1B: out_o=32'b0000_1000_0000_0000_0000_0000_0000_0000;
		5'h1C: out_o=32'b0001_0000_0000_0000_0000_0000_0000_0000;
		5'h1D: out_o=32'b0010_0000_0000_0000_0000_0000_0000_0000;
		5'h1E: out_o=32'b0100_0000_0000_0000_0000_0000_0000_0000;
		5'h1F: out_o=32'b1000_0000_0000_0000_0000_0000_0000_0000;
	endcase
end
endmodule
